-----------------------------------------------------
-- By Jonathan Telfort & James Tang
-- Email: telfort.jonathan@mail.mcgill.ca 
-- Email: guokai.tang@mail.mcgill.ca
-- This is a decoder which decodes a binary number
-- into its decimal value to be displayed on a 7-segment display
-- The bit are ordered according to the following diagram  
-----------------------------------------------------

-- Import necessary libraries
library ieee;
use ieee.std_logic_1164.all;

-- declare entity
entity seven_segment_decoder is
	Port (
		number		: in std_logic_vector (3 downto 0); -- value of counter
		segments	: out std_logic_vector (6 downto 0) -- pattern to be shown on 7-segment display
		);
end seven_segment_decoder;

architecture behavior of seven_segment_decoder is
begin
	-- The arguments for process are a sensitivity list
	-- The process will wake up when one of these values
	-- change. In this case, it is only the input number
	process(number)
	begin
		case number is
			when "0000" => segments <= "1000000";
			when "0001" => segments <= "1111001";
			when "0010" => segments <= "0100100";
			when "0011" => segments <= "0110000";
			when "0100" => segments <= "0011001";
			when "0101" => segments <= "0010010";
			when "0110" => segments <= "0000010";
			when "0111" => segments <= "1111000";
			when "1000" => segments <= "0000000";
			when "1001" => segments <= "0010000";
			when others => segments <= "1010101";
		end case;
	end process;

end behavior;


